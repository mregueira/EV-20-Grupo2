// Verilog test fixture created from schematic C:\Users\Ariel\Documents\GitHub\EV-20-Grupo2\Ari-pc-incremento\pc-increment\test_increment.sch - Tue Jun 02 01:15:03 2020

`timescale 1ns / 1ps

module test_increment_test_increment_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   test_increment UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
